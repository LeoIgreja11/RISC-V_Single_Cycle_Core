`include "PC.v"
`include "Instruction_Memory.v"
`include "Register_File.v"
`include "Sign_Extend.v"
`include "ALU.v"
`include "Control_Unit_Top.v"
`include "Data_Memory.v"
`include "PC_Adder.v"
`include "Mux.v"
`include "Branch_Sign.v"
`include "Branch_Adder.v"

module Single_Cycle_Top (clk,rst);

    input clk,rst;

    wire[31:0] PC_Top,RD_Instr,RD1_Top,Imm_Ext_Top,ALUResult,ReadData,PCPlus4,RD2_Top,SrcB,Result,PC_Next,PCBranch;
    wire RegWrite, MemWrite,ALUSrc,ResultSrc,Branch,PCSrc,Zero;
    wire [1:0] ImmSrc;
    wire [2:0] ALUControl_Top;

    PC_Module PC(
        .clk(clk),
        .rst(rst),
        .PC(PC_Top),
        .PC_NEXT(PC_Next)
    );

    PC_Adder PC_Adder(
        .a(PC_Top),
        .b(32'd4),
        .c(PCPlus4)
    );   

    Mux Mux_PC_Branch(
        .a(PCPlus4),
        .b(PCBranch),
        .s(PCSrc), 
        .c(PC_Next)
    );

    Instruction_Memory Instruction_Memory(
        .rst(rst),
        .A(PC_Top),
        .RD(RD_Instr)
    );

    Register_File Register_File(
        .clk(clk),
        .rst(rst),
        .WE3(RegWrite),
        .WD3(Result),
        .A1(RD_Instr[19:15]),
        .A2(RD_Instr[24:20]),
        .A3(RD_Instr[11:7]),
        .RD1(RD1_Top),
        .RD2(RD2_Top)
    );
   
    Sign_Extend Sign_Extend(
        .In(RD_Instr),
        .ImmSrc(ImmSrc),
        .Imm_Ext(Imm_Ext_Top)
    );

    Mux Mux_Register_to_ALU(
        .a(RD2_Top),
        .b(Imm_Ext_Top),
        .s(ALUSrc),
        .c(SrcB)
    );

    ALU ALU(
        .A(RD1_Top),
        .B(SrcB),
        .Result(ALUResult),
        .ALUControl(ALUControl_Top),
        .Zero(Zero),
        .Carry(),
        .Negative(),
        .OverFlow()
    );

    Control_Unit_Top Control_Unit_Top(
        .Op(RD_Instr[6:0]),
        .RegWrite(RegWrite),
        .ImmSrc(ImmSrc),
        .ALUSrc(ALUSrc),
        .MemWrite(MemWrite),
        .ResultSrc(ResultSrc),
        .Branch(Branch),
        .funct3(RD_Instr[14:12]),
        .funct7(RD_Instr[31:25]),
        .ALUControl(ALUControl_Top)
    );

    Data_Memory Data_Memory(
        .A(ALUResult),
        .WD(RD2_Top),
        .clk(clk),
        .rst(rst),
        .WE(MemWrite),
        .RD(ReadData)
    );

    Mux Mux_DataMemory_to_Register(
        .a(ALUResult),
        .b(ReadData),
        .s(ResultSrc),
        .c(Result)
    );

    Branch_Sign Branch_Sign(
        .Branch(Branch),
        .Zero(Zero),
        .PCSrc(PCSrc)
    );

   Branch_Adder Branch_Adder(
        .PC_Top(PC_Top),
        .SignImm({Imm_Ext_Top[30:0],1'b0}),
        .PCBranch(PCBranch)
    );

 

endmodule